XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��4\O$��ZyZ�C��o�y��������.4s��S��-DW{�RĬ��@����s�j9C�������2����g�CzH�=x����q*��C �E�>&�_�P@.�����+��q�Q�.�Ӄ��S��|�O!i��hoX;!
1HUo�*Ē�)H��c�=����$���5�D�*N�?�	.݄~� �{a���(���� �NYj]Ae@ͷ��o�𼋄�E`����h`��	�	��a�~���ZX�[F,�E��#��%���E�G�H���1q�����'0�$0����e0�����ә�:����ym�aҐi���B��.X��1MUhBn�f��)�-��jT�'G'v�L]����]�����/r��Tqaԏ[gjJ��B����`&���I�Iʥ2-�^�,�̮1�^�4Z�p�M"S�\�{+���ݔ������G �_2dʳS�P��}U�k����B8�����ӟ^ǳ�0�򣬃h���Y�(ySMہ3W��VrD:���������i�m���+t���h�� ���c�b:��>�j��(jiix�m#		ʦ*0:�+�CSHD}{Ϣ:�E3�QK� -|��;M��I}�nIկ1g"��I�Y�~m��%w�]/ȫ��\)4��S����b���Y���]N/ݱ��`�|�B�l�zU�8U;B���8
�B�JHڐIybx���,0�ߐ~XuLؽ��L�VZ�=K��&^�ӽ�`�D|��[�T�of1��`!���dO� XlxVHYEB    56d2    12a0���D���ɞٞKf�<� I��s�z����t��ͽ������[]��î�x��-P�'���p2<#�h�2�vy��K�ݭ��Q�67�t�U�0N�Ȯ�Q�ϊ��.����cmfh��M���T�=�E���yg_�)�̖TS���bs�۟Պ�Zـ��,�����9޴���f�VXg�x�K�RK��{���{w�v�t��<ǆ��
�V����xm�ހ��9�K�b�%3
0{���o:,����_�Ā^ S�ܛ��x�����x�4|�A�<IT=����8�;k�'���2�K�J�*w�utj�9������l��:��9�]
#�9�@Nz�{��PB�(��� ln%����%���\ўp*���uL:@�O\�gb��{�s6m��U�{�{��2tx��������k&I��s�sB���gf�/�����ُ?��5Y&K i�̆���Yܽ1�[o��%����Ju� V@UY!���(o;����-D�ol�v�"H����9��?*VU��!hf ��s �`Ę%�}`��_��@`��3�`�I�i�=l.��0��ͯ���* �����������_��Geʽ��I�&���@����}+���%��־���@�sO#�5<e�hh�������w3m�v��Gvu��W�4�����c�q��;0+xM d*f����U���Hfc�<Y8+�r�扟�������>�~���=�<���*��u\k�tE�DMF��R���-inZ�Pk� ���h4�����,���*���a0ܜ��V �}�^Dt�7a��H �.;ٍc�+̄myw����ߚS�r�
�	4ʆ��!,c���X�o�p,�>���zKB>��W_hv+#=��pQ��]L�	�%����H澀�t�]n��Y*ܟ��aS�F��$t�H�ZD�Fz����I^=f�J-� ��(�\�׮�=�.K%��4?��Jp�z����$t$��P�V]/��ô�����\1]�(͞%�Ў��-��b�Me�����9w]�!=��n�M��̊�")?hQ���_�k���ePJ#MJhNX��/�]�|�D�{�d�������񓪰"�Mc��WCvq�/��B�#�?콮��1���|��c0b�@c�y=���i����{�	�v
���B�r��J��b�-�K�����U
����x�_��~��01�ơ��`̝��_$��B�T[���Bȝ���Ǜ/� ��Z��G�g��.b�����8/�Va�	ũ�ɸ��0u:���>�T}aJ4;G����Y_�G,f�Em���F��r��	�|Z������vqQV��r4����dZW�j���P��[)skO%�\"M|��/r�B50�)O�OR��l�7��1}�9�b��~S&��NMl�?~�{lgN�ʿ�
�%/>SIy���o��|F����wd��2p��F�;pf++�q��&��u�XA�0_�h���R������b�g���x�3��<��}��C��j��D��i��1��Z+)j9;7�0���϶�Nr-N�3�ؽl�BD�A<d	rF"��ڠЕ�v�-s#Ĩ��D�|X6՘�I���.�9���b��!h@��\v�S��i��r��x��ԡ�S}�����R��Vk���>��?�^F&�6�@6H���!ϗ_��aE&����8a�КJ�S������ʹo�4I��6�DE�&	��H��B�����<��Z�k�ߋj�w���#:0�'/���[P*�DO���B��0�n�c�<	�9�N�r�����+-�5�_�N�/m<li��b~��!x�uIe^���M��/���3j�Q4�ԓ�V�^����^���<r+e	������� �Jקc٪f�B���'t[MD��axAp<��?��Q�#� -$���iXQ��{ȱpʄ����O��r��R�9�F(�p����<�(�A�����l�?"x�̟�2z�Wy>��A{��G�4mi=JږK�����[f�@c��Lp}�ƹɮ� �ȅc4ev��M���H8o-�)K��x��Co�s�t��7���ZP �o�ggfD*53�PSkc���C	�L��P�
��h��3?�n㆘#O=({aj��{��]��N���~c��4u�ۣ�s��[�绎Y_�nB�[�`6Jm�̬��R櫇Ӯ���X��'*����ۂ?W��.t���m�K����|�6�>X�X}~�PM�a�I�Ε�QJ1>kxI��O��ፑ`y��� ּ��:`�>�V ٤�@�;&��ڝbG��j�D�����UX?i$�S�
d2��z�z���Y���T�m�{A�� Y=���G�C^��K,?3�p��y���j#�2�TdLxWI뒇K�^����Z���Ij���/D,Ȼ\��2"2��e�wx���%V���094p�/�ĸ(��=���&���$hhST��]�|����E�[�q�%������2� ��B4���RH��4�ܒ�6;=>Wm#qB:�6%�v�e�xh���TW�A8x	��6VR.K����GeBy_q���
�se�JsN3��{��hd����I2�������4\����:��L�S��U5t0�b����mX)ĩ��v����(���N.����� �zLRD=������#>��:�TĒ`ц|����)�_ݷ���|�	NYr,�i=�wp�7�K��Ք58�#�����J}ŗn�_�T����P��I�JoB��?�?�K-�&\�N@�9�%l,��\LΩc�$����l����0,A|}�cW	W`����Ꜿ�`�r�|��S͠H���!��Hn��3��+�s���R���9E���.�~��0'��.��X�m���^R�y!{#�4o��}A@з^n�j�u��r�G���� o�ڮ�+�SPo7�W�gva��l5��L_=�)b��l$�>+�"D�ӕ��,ɍƟH�#�)w�<tF��c6#�|����f�|�Ӝi��~�?�mN<l=t�qy�ڀ�T79Kl,�L����}�Sz��߈�U��B4�9�@t������t���qNZ�d�6�*-��e���tE|]͟��{�%���D�a�D���ii���=�� �ݷ���T��7d�C��Ь��8�O%��F���C���".%?�u!��7���p�?���c�������X����.��b��^dc�����'����x�P�`�F~��g�����O4�HB���nk͠P�H��D>����p�r+Z#�����s��0R�I�-�X�S_��P)�����:-�NJ�=�-T��ݾ�b��?)�@�����I��y��#���[��6ш�\q�c���� 0��dWA���'_��+�ݛ
��r�l�8%=�בz�k0�IrD�P�pD�����N�[#��������L>g��Ϊ]��m��	Q�P�<q;#S�ϱ+��˂+nm �p+��W�!?)7\w^O�V�a����q���䰈Vߵ^+1k�_JT���f""T]o�+`�"�z�mG�`XXp��ښ��ľ떃!���v���S>u�ǁig���*~e~x�Ӵ��#~�$q@Q�U�$��֟�ecO����t(�܃�R<N^�.��m�a������I-HP�0��u!���a����e��b�~d�]�V��gld#L�U��[�e_F��0x&��ˡ���2~��c  	�[l)����vW7�����߅���<�MnuyC+L,�hMz�Dҕ8���tk_�n$���i�JKԛ��°%2U����W�T����L�po�J$#�'����$ ���*�úL��:���5��pp�Ĕ�������$)�=���}~`~�c���J�}_�dC]X�ȍ�e�s���U$�����%O��軇f~�q8��9HDv%���F}���U���>��b($���ӎ�⽶���mВ�n�Z3�ٯ �g� ��(���#������������	�{���Դ��⓺AV�#��R�ֿ���n�����'�/ס��c�> y1/�؀�f�-�E]"	q���Ē��0���F��D?�D���l;�r3�4��BEgf�}���?g҆xO)�sG7.���[���t��}!�w���b� ��N���5�E�c�Bv��9���
�+��1����g�o�o\+�S�^ �2N/��ɇ���x�S��w��qsąǳ�����R��)�3i�޼t�Di���}q��A�Ɓ�� 8��|���Ÿ��+)����k�ʫা�:@[��֢Ui�n�ߓ�9�" e����8���/B�&@*IF�]��ޥ�>�͡��A��sa��j���wJ���F\���vؐjNt��,pK��-gQC���Q�O�!�~����n���_�jכqӵ��B��v��� ��M|�E�A|�_��>�2�;n��Y��	T�[�xo���zZ�`a��V�]P���t����U��	q�g��S��RDm<C�~�R8`{�TII�*h�U�E�l⪪A��	<=5
K`��9'�B�,)��x�3ۍβX��p�_G��P,=�0=.tY��1/&_ơ�y�^<8��B�MV<@$�*/��|t#�p�zD�ȸ\�s�V�~&Q���v2iƛ�fSx�6wG�#*�F