XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���o�^�W��7��mp�b�ꚰD��o6G�l@J����E�e��\�kv�O�	����.��|R�CPL ���P�4}�Q��ԅPt��И���i_��/ؠ9�Fbx丐*?&S�B�������
�g�O ��udN���S&e�]c\R
0m߅6���RA��E���^dQ4zr�x�L�k�U��S拓br	�����y��سU���g�O!���>���_���&2�5�z[Ưdw���x�p=��>�$;����_dgntN]+P���P�!��^{�J�w���2���Q]�@G���|DEӁ��!0�~����p��f�(V~�۷��C[^������>n�]`{�o�rf��,˼�譀z�c��s���$<C��Հ'�躠1g������ig�e�o��-�����@��-�..Ht6d
Ҩ���g�B��L"W
]�l� S��H�c��b�a��M���%A���Û����5|M���/�9
�h��	��4ś������ÚC#�f���ΉV��P�t&E��%�u�.����a�X�[�I_��Kt�[j�]bE0ٷ@ \d3�Ϡʻ��z��X�U��Ga��1���[hmK��-ށ܂a��wW���� X��������Q$�D�|,�c5Eⴚ���{Qӗ�`$p>s�����$=̑�ܥϗ�+����A��B
�!�#x��z��t��P0Љ>2�a��t�e�K�5S�:�x>a��Bۯ�uA&�u�G�^�@�����tAt�XlxVHYEB    fa00    2910���MB�?d�+�Q"%5�-:��+�Dv֞����(�����\?����[bޅH���+����Q)F��T��=}S��5��p�7�N
d��B@ ���Zc�0��/�V�`�Emc3u���p6�L�� X��׎BM���7[�ڮ;F��
���W�ިU �ڂ(��i��S{�e�&��0wkP��-ub�G�;�b�d��u�?�L�S�ZB,�XGy�Uy�[�Yz9�����鯑�3�_��]��هS_���_N�w��;Dփ,�#�)d���z\�ŗ��\{�yq.���
�D�� )�-����S>WʏMŁ1�Hԫ!�2�3���<o��}���_�Ұ�������g�إvf��B�e�o���̞C7�Zc▝34}�&���3�_W�a+��_�9ٜj�B��x�!�/<:�g1�f�@���F���)�_<aѠN�"S�t=��j>x�2ђ�Fh�-�l_���)�sR,���"GU[�r���N� �6�{]�ݗ8Z0Y#k<a4L���;J�G8�p�wý�H��X��T5-��c��u-c`&�-���g�W�S?��4����]��Q�s��u#K��U���N�����m���f��"Pf�N1�	$��?Difp+�U�����ة���W5B��~��O�(;�(�d�����OX���<B<ʟO�Cg��	�s���26;���?�����zf����DĸO�1Hyg�#��- ���o�i;��C9��)��a�r����o���~�1�uyM9�6W��/h��H�?�c9(�ٱ^ _���yL4q���(�v&�a$����[%Oa�l���1���K��̲ч.Ԅ�H����/��}�&����h�I�K�WI5?pe�^9ژaZ9`JF�f�٪Q=_CR�,Ε�HFSK���;��$�K��`>����됝뭜�T2�qH�j�k�BoSЯ;�wg`!�ˈK/���L��d�d���P�B^d4�!����=���A�J;�Ǘ#�bĚ��L^���OTg>�Jc~�{�0B"�p��4�n��k}Ns}=G�r�͉�XL�M�:�覾�&���5��bI"��\bo��'Nǩ�F�#j`����դ�G���X�	%:,��zwO>�6����"�n����PJ�h������[��f��'Q����6�ڔ������)�eU���K�]�Ǫd�z��	�#i3��+[�K}�D����C}e<�c,�?9�����eih1��	��L�<	��@8�y{��Tɗ�<m���Ze)B��'Ւ�e x7H"tJ���Q���o��TJ��FNf�js��aᕕ^'��~�1��@�؄��E �5�1:���7)�Ȣ��m�w5�`�DP ��@�DD̑pv���x���ߚ']|�)6(�"�h���h�tW�'l�W)��Y"����S�flI]��䖧�q�U������iLU끁'H@��ޞ�&?Wq��dÕ�uP9��$�d�B\~�w&�9箬_�g�����+]�9�asG�V�-8�pz�?lQ�_U�eB�i���W'|�=+�U�1բ�M��L}^���z��8��^-��|y#+����c���G�ZF���-I)z���m���v��pd����H]�f�\�ɒ~�)?�2Tڶ5�,����Do�\\�zw���y^6, �^Xԥ��u:mU\K�߭'jK��1Ac�u����΋���[]��'��uKey�Vǈ����HÏZ	�Dt[o-����2���[��v�*h���R��wf;�JA��?X��j&�� EG^V�t��5��
���7�>�_��ܝ�'~�[�y��Z!���g���񬾺��s�kn.��ܒ�b]}-L��	��^3������2��Js�qy����c��"���gGNwXh���32O���:5H� Ř�ŷ��Ԗ�冏z���"��s�bU���QLÅ8�+�MG�9���̇ ��i:3��G���Hڐ��Q/��b�@^N3Y���#�yr�<�0�sUP�Gj��׀^��c<}�r�y+��ه�^\lO���V*`B���ѳCrK�[R �����φt/�ҭ�Z
������*�kU���6�D͹��n[�59�sT�^M���y`BI��?p��
Z� ��Qr������
����B��]}kSVDbŰ�x�D�vd"B����c����<6p��X3�}�WX>z� (�@��������ˎ<�S�OD��( �s�����k�C9~5��R�)M��qAh�e�W�g��bw0<���'���^D�h`��~��?1�a�5;�1p�Nb�EX��y��[q��>��RъS����Z�%Y�wG�E���� 3|R�[>!��t8���#�h��׍A����(\>�b�ek���;�ތ��0�xs
_!��*)�X��Z#�k���A�Us8:\�̲�%��I������~�B�ͣOTo���9�㣮#�"J�I0�=\!�u���i�A���(�^���ОS���Y#���Y�s�!z4�}~�_Ds�p��*�/��4l��x,=�Ɵ3��h 6R��Z#�9�E-���M��
s���Z�"_u}�|��r�;�2gg�����0ב��^�՚e�"�3��A:˼�<wJQ[3�2d����m	h��ƀ������9h���Н�M'�c�v��0h�6:G{�02���J�s�d[P*����Z'��0Ä�:���n ��G�9e��y� mV�w���ۣsyJ2)U�[$NWt7c�x�P\.xV3
��\��?��T�-/�8\�$&�+2h8�m��W���:@����o��y����b�4l]��6�2h?�"w"ZN{@����h��n�4�|�|�9;"$���|\on�>��' ��8	�2�-�`�h�9�}s!��v���n�J�R�3�� r�	>#YR+�''��)��oY���C#�����n�-�9��c���nU�E�(o�vIt �_�˞z���ʄ�o����p��B�6��h�y�Зo"F� �k�+����p�O�jc�~��\ob�9�$�ʹڒ	m��[�������U�{j��_��?�+�SԄ
�l��7Աu��_�X�5�Q�!�G��(8���]�5�M;�dexn4>��0�\}��J��<t�X�T�/�;��(��+�Kx��qH��t�7�:�pq�=b���!�H�~�a
�ܳ���#����p��:9� Jh7��cpﻦ���E��pGBѲy��#D�c��FlW3�۲a:�ڴ��U:��c�h��r����%�I���&�bJu���E}�?m����� �E��T�xD60�!��b%��߭���Op.�E�����V���.����~��q��r&C��a���JFs*؞�=��T��1��^sdjy��|��A�g�[}��rw�OH�`Va�rG�'�%�� �nLO"J �4�{��3�I.�;F<!���l�gD�j�)�47?����l�&[�G��cj=fHkSwF]BV�O��J�o��X^��d��))tЮY�#�4������֫cI{��]��ӛ,Hz�!q_+�⤶ޫ���<A����7�������T%��J_�I�#Ȩ�c��[�8�:V�vPz��"��sȸ<�c�S(������XZڀk�S��i��0��
rF+�6W
nA��F����"�b��F"*�Q�g)�0b:cl&h*�6Q8�?� ��*_d��V�44�[@E��ˡu���3�)x�Mi$��I�B�}q��D�(,P����Kj���,�$:o܎QV�n?�k�R$�v��~�g�G�x���:Ӳ�=����DfCA0.��S��q�u�t��	G�`I_[&�7'�~E���k�����zIB��x�eU�ɶ�"�@���b�%�ٽd���Ol{�GF����v�y%oS��D+���Q# �^r%ģ�?�v�X�E��/b����Det<�[�k�����=��`Gp���͸+0����iY������8@M�;F�o��lZ��IA��������G��D�y���)&Șt;�u��l��4[]К"���C�c۰x`�Z�~Kn��O�c:B��^+"�?¥�}])"�/z޲��'N��[�+Ƴ
m�T ��5�����-&����r��J���	`��Y0�(�m|�9�ltTL5}�ڊv f�p����Y\.�m��7�Uc\f&�Џ��0��=�e��З�l�V��C��a��;JYMњ0w;t,����1L��=�V�S;�ѡ��o�Q)Љ��
�x<uR+{K}4�V��C�H���/���:�Xl]�>hMj�p��6�8~���.�<�9����׵�SWl\���fAe���mfp ��j����c����CarB5Gv;u�kW��,����	w�Vg*�f�!�1l���WϕQo�[����rI�W	����&QbB=׸_
��G{�<5�xo�;(2� �?��Ԡo�\s˅,ᎁ ��EPZ��q1g��˦6�2��}
�[v�U���o��L_��x [�=�
C�5���ވ��d+OZ(��Ϥ�Ԯ�g�EHPt�C�%��4�>#u�7L|p����bI �w������V�G�K��'X�����3�ψ�Yi�c�酑?F���W�48�[�\xE�|����SƯ�3��|������+�(/1��6S[�>�C��P���S�,� ��}w�p[)�M7z#ݫ�GvI	�ʆ����Sx|RB���UW_������;��a��J�yS��)�0B�-i��F\��q�{���23A2�m��ɛ �-���k⤢���&X}�6�f����č0[,9�E�k�|1�4����o����R�����'~�%ս~�r�Ql�������c<����4�Dm�
Σ����B���2"�ZUD1�Ϛc)���=�ݡ�%I��>eu�����;37�^�t� ���"X|V��2^�NYIr/�iϣ����$s�X��o�F�\B~��Z3ZX��{�9ekC&���(�4�F��Zcs'�k��+�����=|@��XPK�F��Ld �&؁��c������B�p�h����N�A6�f���2��犆@�+;rN<R2���4m�&�z4\��^x�{}���t�7qrɲ�8�!�T��Y�t����F���>�s�~?��V36LA?m!o= �U���*�C���E~S<,�.��Oc�/����xs&�aq�j1xy�i��n�޻�C)�Y�mZV@ρL��=��V��R@�Km,�K[�ލ�*���]:�F�c��=�e�63ۤ�A|��Kא�eI.l�4	P����v��-׈�i��+�'p���H�Nu"y~>��Q�D%�[yx�iu��݀��H'v��b�o	� �����m�D�M����% ���0�
�ʻ�@4ģB�\�1�]�-��
�p	�6V�i'�h<d���S�bh�U��ˇ/�^d�in���<�f��G2*4�Rp?� �:���(.ƝY=���sy���Z8U�Wǝ�� ~y<S����Tl�8�/rs�t�������]�=�R��
��=�HwJ�� J{�[��%i�=�t��xi�_�o2[�g���S�P:��RZ{ǇN!�a�k�M'��j.B~�%�y;I�iG�[��+)��(�/�$q�Y�Q���ֺ9O�S�٬����6˾�L�`x�"`��<G�`"�f��fǦ�.U�S����#�t^�?D\
�.q��?4xj�����5?��9�s�Gn�u<�+���LB����+�s�؊�XW<U�AG����@+���FVol|��^�X����H��IK��v���qj?���t��58[�d?�xQ��
2
g�l�8Ͷ�ʡNC:C��Xb�`�ɸ�0c(a#	=_����|����Ph�����A}[�Ĝ*�,r��q����1��IvS��?WFu�Rru۰��9jP���v�,hF�WY�"h����R٨e����FS��.����OA�k5R�xح{��@�"��S׀�"����b�)K9Ӓ­^^H"�Z��3s�tq0�����9����oc\��۸D��h�b)`�~�:� ��P 7ЂMO��*߅"�+}�ɛ����up�^)��á4�qL
�Fx��u��T����>��c�J�ط����׆�i[���EL�B\���X	3��؂t�j�f�w���3��1-��@��ml)f����k���K):��KN䦲�T�>���W�݀��a	<� ��\��w�]%�U��^�8`SOP�َ(�{��+`t�y���0��z�)�v�3fX$D���N�ㆶ�8&aڹ�\H��Hݛ����\�����lJ8�����j�i7<Z��=�����ˀtԍ{%%�Q��؛n�X��{�HQ^,qg�'�|=�/���z�Ε����jMƾ8q)��~��g��uQ`���v��
��x�$Ks,����z�wm�DM�w�C"6�ΟŪCjv��,���~�u����1������J^������T6�B��iE�)����u��Z�kl
-��"u����\�H����w`y��a+w��#�U��	{���V�"�½>=�[��J�qꮭ��y4na�����x��[���6�H�VhIa�J��S�y�>���+x�Yq?�y_6)⁛�
���מ��A��/���x�$jjgɞ[����5�c��w�j =� _��v��������^a�JT۲E�(T'�n
�9Gy�LW~��m�q����*�&v�*DKZ� ������'�ڡ�X�`7���`w�un��y��v_�/�Fي��օp3�����y)Yt���p�X�{�q� ��Zi-ai�ͽ���`� 5i����]y��=�]Ej�C���Ѿ%?�U�чn��K���دˈ��ht0tr)��H���9̽>����J��j^7�p�:ʤ>��.1˶Ϣ�.i��U1�����mH �n��2 ұYA��k�_2��,��Nu���a�V�p��x��z�K'���N��s�&���������+O���4c(��/�y����(��I�~]8H�$Z�U���+ߌ)�W���{�`hD�a�ꍘh{�|0�fcԬ��%�\!�N`��4��vM�l7���ؼ��zmZ��"�\;cp�Ӿ�_�`_�ߒ��ٰT��-�OEFaW�sȋ��;���V]d��\9�Ob��65R��z��9ԇT��"�;W<&�Oz��?+`�Ef��p���3�]�H�+;�Ai�P�:3rK�|I��NJ�Sb1�� ��W�-`���u���f���p+��� &DP2�Ol��yֲ�m+���S�EZ�=� @#�D�a5����2&���z��v�v��5���%��@�Z!�K��$��	�1�-���OȊ+�f�[q5_e�yH���\� �9�T���������W�O����ݘY4ӵ�3�w��-	����*��A鼫6�ci�=�L^�vKFT�Z�ټx��8����:�3~��e��{=���
(�ۈ���J"P�̻�m �?�q�y��G'��M]a��� S�5��g��X�Ȧw!�$wv�-�hL�F��v�+����w�L�S	j���A��W�0��� G����+�R��Q[��Ý��+�8�T~.��6��&IK�#�u��\�;��I���I.��awg��KE�W*CzV[p�7�Z�F�jr��io�ӆ,�e�*�h�!�ȯ�x	�� �b���ʭ���v���$��f
� YIa:`#�e�֋�w-t[	�����J�Y|��z��"��_.���2�=>�hm�\9[/c7h��<l�����R���jp�nݸZo\��� �T��Ղ>����Cª]1����Nk���`��嵸ιŶ���@���FND����k��inT+��uġ����Bn,L�t�*��_ ��$��5�X�_ҝ�*,@B�q�iQ����}�
H�T�E��/C
���lX3W��,�؝�5`�<~.%�Do��<ͱ!���1w���=꽇��H�;�m��f y۬��#D�٨H�i�Ϗ6�a�78S�#��nE��vB��O�x��Næ٫x����f���P�i���rC�����Ψ�P���*�%��[1�ż��kT���@�1�Cn�8�,��4Wč=�_{�A;�b8��c�Zc�Qb�)�돧2fبC�,�C4kD�\W��:,��c���@q�M��iiH�v�+Aż��"��W�C*�ќ_�o�TR8����+M�ݓؚ�H��N%� �>~�i��H�F��D*��mĳ�-J�"@ޙ$�^�IVf�e��$w���a��H�m�w��H,����u�9fYS����ɥ
�ٰ�&�w��b@�Q7[4�Ԇ
3먁]٪���P,Ps2;�
�`9j����N����G5%��
�[
�;��@�e����AD�}&����>\U5-��-���;�vE"TY�$ }�b�R뢉	{�Rw����>c^��FU6����Vc�����n�h%$�Hd�����؈N0��M�H%Ar&��T�$s̡$�;��.z��D���M-Ii1�M��C�XAzU�TB��iyI��T��-�[=zg%NaH����7\%��Q�>-B�̼@('�הۂKɨ��q�çIZ̕	�5�|H[<�Y.�,}�ushD��bi��U��$ �$f�I[����
3k�2͔H�a�a�ܤ"���a5w����p�<�K;�%6�9�Ts��v$J���Z��0���=��ڽ���h�U�m�����m�W:�>���ڈ���I�3]Fz�H��������H���s���&@������f��Eg����N"C������Q�H���� 5���2�}P�0��� 'C��=�bg0���0�����a]��>��TaɊ]�p��A}��o�t��~�w�!�V˛�D4�:�s��W)��1�O×�$��n�2��`S���������X�:��a����c�م�n���f�{���-`������{�WEo�ъ�x��B�7p9:�Ǧ`��y	�7���.ic0��{IZ�ۯe:-�o�R���o�d3\��I`��`�u�hzUr�V(wIKN��k�޾�F	���3��y4�;3�\޼}��:Nnd��s�a�ٗ��N��p�D�Z�#�2�ۜ���lg�Sq��:��8�����f"�n=��B��J[pG5�97,sy{Ӕ_�����[E/[�,*���VG��zq�"U�������`��yKH\�f)��Q63�'V)c�&O�� {���'ܪ"����\j�M &ɫ�G������|��P�?�h��7,zh��"��&L1�a ��������2��'�Xo:�W�r�[����o5l���q����U]L��uR�Â3������J��B�3�~����ȏ����=�F~��Ḩ�N���ߎ�]+�\*I��3�W�J(ZlE�M,�ix/L	�5E�?��Jp'�
� ؚ'!i��KN��)�C�}/�T� o�,�e����W�-�0�[�?�>�����ϒ�|��@�_ڸ �?Fv���U�8LEX���ZBCv�xφ�h���"vJ@�eଊ��Η��Q�2L}�XSrߐ&=�C0�'��2z��큵���n�/�z�
O�+�����i޲B�Vּ��4ud�b�����)���a!I}��GŴ��{�n��ς��Q���&IKnN�F��4���v�~�|$o}�����.#%Bѝ�?�1��%<d�`�4�.�>����qB[79�\���z� zy=*4i��n����W����X���fD_Ǌ�K��k��O������Z�{W��mJp���Dl\|��I���S��Λ�0i�!�	�B�	P�>E��9�`�A�ڐܴ��[��e+z�ZTW��������E\�F]��b���v��'��w�F����Ξ �t��32Z0șWC5.(e����@7V�%0nk��rMkK�ιX9o���O�P�~�!1\���5X{�oA�ȳV[��O�����~�Lx�ꀚ��h�O�+�-�c&Fh-.l��%K��8~��l'��1N^&��:L�ݐ�8��!�;*`�2���_�}���˻b������O�kғ���/��e,��Mh!薆v�O��&�?��4��_�
n*��֞M�-�$O�5 cr�F=��4c 4���L���A՛ج+�TOvu�}`��Q	��9�\�*��w��lpk��?h�����B��s�"c��R8�L����Ft��{��:1B�~p��pw�L^;yXlxVHYEB    6184     f80�|�*3š`Q����k/C	�@;P�*����q�ܺ5MS�D-�������Ym�I�/b|�P��6s���l��A(pm+Y�@���G�I�7�>�w|Ԅ�5l�c��+;�DCE}�R5��BrHŞ�d�tt�~��cS�:݋AYĈF"O��'Q��e[��$,���L��u8T^M�1��)F��t�;N���ظy���g����������q�~�Z��:������������t��_7}�r%Q�O��+	t.׽q�Ωb9��O3>��H�ǽ�	Q�7����������2~Y�H���nh�~~
Kl%3���	�GV/�o+��w�Ԥg��3o2K]O5���٫^�LZ�Ú�9yYQ�J���Ǳs���bJ�=6�l�TK��ک�?��.|��Q n�l.������!�@X�cUJM��jkjm���]#�t��l�b�vw�˼�Ύ�ӂκ3	DNQ�Rƚ�(�,�������)�_������\�[[�x�����չ3���Tv���LH[�q^k'�JÏ�V*�'��Ϣ�\�C�"Q�;� cG�9+��T��j��q�O���(�cWp0��� O�eT�� 3!XΙ���5����� ����-�g�����B�%N}*��1s���EPD~��עX��A>Y��\p�Ԛ4W��Y8�N ���G噿���s����,:�e��#MfK�gu�Y�����\�GY����|O�rτ��bl����� �����0I�HsВh3�]���%b{�ϱl���k6�O�H/���n���r=\��Q�����+M��7�LW�Q>۰�ü����#�JZ.w�����8�__i
��w,��2��d��R�;�\f̀��N�_�m�%�J�*NM���e��l��q���٩�� ��",�wk��J�N�2�_�)� �ٜ5�'ZSo��C�i���������
�Z�3t�\tY&��m�W����@4.�) g���~�=�*&�#b�iy7n�� �QЯH�yp�+��,S<W%xW'�gP�e�:[�*��dd���I�"�v9��y:��f�q�\�l^�@���3e0&֕���?�H�v=1����+O=:�0[Y����)��`�M}�8�/��2֨1d���7�]���H`7�nfA��t����ڵH��A�D{r�a�z�PM٪y&S�.�[2χ�#�MN&����z`���_�^���RUH)�"-�O��� �Uܢ C�̻���iQn�Q`�8��l�1=����@K�� Q{.r�%`;G�&����������IF鯮g��cQ��S�����*�[��v0�b�R5lX���ڵ�]9�1p�l��y��Lq3yt����w%�E�WF���:a\��]��vC����i)�$y�DZ��6w��9'��#,~q��2Emw�ޥFW:�<o��	�D�=r�\E�}��񮄓�MRj��´6@؆s�[���H"�@붱E15����7�I~�0�SX��i5h�������d��Q�K�@k�b��:;�o��yM�No@2��P���Ra����$Д���0�˷�݉C�l��X����q}]�*�z;R(j+�C"�|g�.Ø���A���|��� ��/5����wjE3G(���W׃i
5ѧ'��^@n���)AFgfǯ�7C��� RjS���}�ΤЅ:���B�֮N���[���'}�a��F�ѱː'[W�b@���3~fWry�ȳ�fU�AFW����'�j�e��-&�6La��E���� #x�{M�r+F���)�4Y6�(�i������K3���\n/�u{:��P*�
|���Ydѧ�_&}���cG���R�B �F6��$AN��^�Ӌcs�|=/曅�K5:¥�O��ފ]V���7�����Ő
��r�3����A��j<��
�oj�Y����*��TWf�~��G%�W��C؞���e&�m� �������p@W?%̯�Y)��d<B5������P���}�D���"萿��*YaN�+δ���M�d0q.�M��P���R���Ɋ�v��LZ!a�?�ߴ��7nY��Q�,�hڳȳ�Ҵ��M]N�*���� �Q�Ӱ��g�J���]Ԏ�����9��,�x�q�:�%[@�k#wo:���([GGI��a�4&T�tP!�W��f�7t�X�`$!þ��	�˛�vg=P�_���ll�+(�%�u.�gy�3u@�a��R�ʽ���=~;�C�ߢ����Xkv�o;��B����' $��#�ܨ_����$��_���hW.,�TĲg�o�Fsj��i��_L��Yju`�	�G��#N�л�Q��?c��4�;l"^7pw�h�9�u�%"��CX���w.Nt��Mm�%MuW�XIu��w";r�� �Q=��4.#t�#~��&{yЄ�k%�a�;櫓<H�֫
��?~�ZQ�$^���������FEb�������u�I��pj�e.[���)	�}3�wᵵ�ɀ�i�W���</w(.��<Ux-�6K]�ů_�2c\srG��Ձ�.�Kn>������针nK"Hܘ7���{$��]������A���l45E�{9����J-��֪��9��?Iɫ ��%�Y�g���m�f�J$�E��8u���+Ipq�t���~e+Ŝ�F2����5@�O��X��J
�	�n�����/3�)�� �#W/S�A���s+ׄԈҞ=���1/^Z,� j����B��?�ڒ�{������$�()�Px�&�Ƭ35
4}��X�	�?oRP��Y�uq$s��Cs��BL�����A
����)'�툺�T3�&�Ȱ��'m���έQ�b�]��i����w��K<��[̐�6�B�K��n�V�Lr���y�KX.��E!� UP������ qa�y1u�ݨAf�[�?��1V�&5pk�SG웯&%�]ŭ�����y".Ezr�߲S�rB�ȯR��E�Y��M߼|��ڦ@�J�����~$�Yn�u�R�w^Ȝ1{�Aѡ��w���3ۈ�$���xa*�U# �C�z?�����~���pF4�{~	!8y���e�
�]�!��]�(�y_��d�� ?Jt֤���.B��a�O�s*�^�a}�7�]i��A�������COo�.E�s2�LX����=ݤ�S�9Wu՞��
�+��Gr� :�]�+<��l��K|K���cBJ��g���Ţ���.}Np�@�uJ,1q�|�x2ma���f��#?>���
Xn���Ig�µ�nD�cJ�W�T�4c��}�n���H^~��A�F�����&��xU���/��Fc��Y V�q���컫��ˇ�H����<4O�62�l�������8Yu�(���9��f��^O�O�dh�=0�Ŧ�/�I���xI�h��&��F1�i�"�����~��l�4�/�����Ipu�3��'nU��p��L���g�h']@����m�*垓�x^m�f�%"n��	>h�#'<�Z��$��4�*��?|��O��d-F$a񁩒��U��]T�tPPKa)�F�Yf)u�r\�#��������A�脺q��\LFΪ��$��W�����$K�ؙ&#�B�m�8��A}�*8C�MY��+OSL໬����HL;.7m�� �|m�P|�gQ�J�F��wү���+u�،~���I��o�`?i�*�6~�Ɉ�G���}��i��������������� j�������^n����i�S�8I:=.l��螦�䈊���'s���pɣo����T<-x��j9��g��NJkf�
�
�7D7�����Q|b���S��]�i��E�_������@Xl��