XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����=�[��@R]��"%d��¾����o4��Zi�\EeD�ɪT6�RՅ�?�f����q��6�y��yh��R�<pZCٸ�Hf��pav�(�V}?B���E��~�=O���e{��x��7��`=J��r��i���J�^�׋��W˫����í| ���q	�"#3SƎ�J�>G%%%�@{]R6��Za��\\���X��������of'�egU�e	���`�a���i��s���:#6�g꽣��]�o�k��-b��HJ!A����mznWr�'L�<�x`�='
̜��q��B{����?}T��,���XzRr\bҾ��1�|FC)bq8������� �Y�1hd��۩׌�$�.���Ղ�8���X	ՀC\؛�`����aU�1��T����?����u`��:�@8�9��M����Ͱ��Pn�A�y�u9�Y:��iV��4�B�]aw�)	�b@���ϳ$۫c;@�ϥ�F������Ŷ��=��Z܌�'V��� �ɷ�\$N،'0�^	,f?��Ic�g�9?���+?�)��K�;�&�j��0�Űo:קZ}����d�!-)T���۫�>�Ar�o��C;ט����E5�e�	ν�+1Y�n�J�K��u�)�Q�(Z1r�L6F���d���p�<�6K��c޲��	�������j���cW_<y��eJļd�A�b���4$�|��!0 "n�����<���P*Aa�u�[��,Dހ�9}��@{��zXlxVHYEB    2e55     b00�*��T*ZT�G �W1���k4�e�*˶�ʮ�
���ȗ�d�ntm��S���&pM�nb)�B0���
a��&Y�EA^sC	r��2b���4H���S������������g��*�l��A�:j
DS�R��'"��̎(�{)	İ�����=m���h��M�,X����{<z��9� _`rӨ�	^4��_��[�엷VC���@&����`���V&r��`�)EĹnF�;p6���SG�7/�iA�LXQ��{�	�����Zf:N,����d�ͱ��JX���Q�?XL��Q6Lhd�.�S֓���BoFŅ��+�D�_���A�۟��3e���z���-����M^�j��%�!c�6�E���qj��J�{�Zvr�c��@9����=;}��J�л�=vNc50��o��Ԡ�ݧA@��('�����xR>�bZ�)�~�����u�b|�e��0���K�|�0wׂe��zS�s[��Ԣ��h=�ϡS����k�Q�ϳ�5�ꭑ�9���%����Qg�OKx'�q;LqP�Aoh�|�����0�M�^4x��\+C�B����W�t��H�WOI�X*/��ˡ}��B�i��f�å:E��TqR1���/�0뼏`#=�|BU�ʨ�03;�?)�5�T�}��"��k�qQ��&m�^�̭:��7�[Bq?5�_���mZ�����4WLu�-	J=N�\i��|���dE���u�+���pD�;n��4q��W����1QYt.��ѝ�~3"�;@t�����P��ڜ!D���
����D�V��n?�o.�Y���bR�S�ͪ��Q�e^����	f|���[
�s9��P|���>T���o������-��>���{���4���/*�ȼ 5s&���Nn�Ӡ�Ua	�$܌��&%��B�P���PK�q1K8
4=�$�~�/0�U�r����dU��:ʪ���������5� �N�Q�KT��5��[b/�n�i@ ���͊�#; �dw$�����j���e�Qq �����e��5�T��蜹���:�ʳ�v��mK:�HL�}�y�����>�� �4},�,���%����˩(�S�7�xM���ە*̯g��#Q,�2	��!J���!R3�~��$�SA3�l��ߡu��-|��Hi�� <~�����`;%|�n����RL��Ea`c�� W�r4�w0l0��� 2x_��â�w��y����lSYBft���\3_�������(�fZ��L��S�e�50l��ɪ^���3��݉�&[���a��fX])�$��A�3�P'�#ʴ�`͢){Ri�����聆���<���z~(�R�4�.9�� �t�҈��9��`"������J�E�f|��1�Y�5�R	SH�@Ja�,��J��"�CN��8� ���T
*�q�R(�h]rK-���Q+VU4t�#�X�q35�
 G������_�S��Aj�q���o���	ƃ�l��M4�e�l#!$�M�7�nQ�"v�fUVŲ�Β���7(�����N{����#�FF���(�7����A��t���h�n%�2w���Y�2~����9�X��:'���8�C��*��%�!!h���Ý*���w󓿄�fQ�Ą�GR;��Z���u���T�	���������:��N�z�r,v� ANn���� @+x�T)��N���S�Y�c��]ժ��{@�[��+*��%:��	�s{-,�[���`�l�ۉt�1L����;�K/������0K�]�CN̬�^�<���(��Tc@����0�$�r�Aⴥ��{�՗fڒ��jO��H'�E	��K�VPTTW�_�|���XB��S��d�?p��p;ES�����-e�ѸY��qvN,��.�����[�L8K��&��{! ��	�3p��T����������>C�/P�DZ��������ᆕʌ3�o����K"�-c��Vc+ɊL��{GdV�F�)��"l�|��
�H���ՄRϏ�
�*I^1��*̕�uo��~^]2߼�/�����L�8���J���i��~Í2<`7��_^�S8g�>S�K�;�Jq���ՔaGr���z��_���[�izB��͛����2W������}�%���wRL�,6>B=k��Y�����p�P.'�T�͑��aX��GH����� ��.q�#�?!x\P�>c���
��ں���;|r�}��zӃ����C������㞗³u����t��"]��:��������:8�3���znt�9e-�5�M���`�p?�`J�"5�H��UZ��row�v*L���!*��R5�t����eD�v�6��(��\�hnOXʥ>��7)|���̡�m6��'���3�sf��t�9�6nAH�"I�0��%���ŏ�n�^I'���� ˕���2�aXVeE&���`pA��Z@����&_�7�y\�t�D�:������� ��┟�O�,���~���O��v��˾h'�z�g�K�.����`+����H(�� Hu���Λt�+���ϼ�����c��=��7��֠��ޝgz
w�"��{�!��j�
�����q���{��\�U���U���tƬ�J�����Y�1@��H�ɩI�N֔e���.�� K3����9K��u)P(豫�O��|]��c�hLY���VӼ�Xn�HxAX��-w�FrR0���_�KL�d\}(&G�K�.���XF��k^ڥ��獔�#�X�Y�sݵ5�x}